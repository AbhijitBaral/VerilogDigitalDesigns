module Exor(input A, B, output ExORG);
   assign ExORG=A^B;
    endmodule
