module universal_register(input data_input, sel, clock, left_in, right_in, output data_out);

wire [3:0] data_input;
wire [1:0] sel;
wire clock;
wire left_in, right_in;

reg [3:0] data_output;

reg[3:0] reg_data;
always @(posedge clock)begin
    case(sel)
        2'b00: reg_data <= reg_data; //retain
        2'b01: reg_data <= {right_in , reg_data[3:1]}; //Right shift
        2'b10: reg_data <= {reg_data[2:0] , left_in}; //Left shift
        2'b11: reg_data <= data_input; //Parallel load
    endcase
end

always @(posedge clock)begin
    data_output <= reg_data;
end

endmodule
