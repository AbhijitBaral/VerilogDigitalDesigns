module Or(input A, B, output OrG);
    assign OrG=A | B;
    endmodule
