module And(input A, B, output AndG);
    assign AndG= A & B;
    endmodule
