module Not(input X, output nX);
   assign nX=~X;
    endmodule
